.title KiCad schematic
Q3 Net-_Q3-Pad1_ GNDD Net-_Q3-Pad3_ BC817
U2 /14V4 /14V4 /14V4 Net-_D1-Pad2_ +12V +12V +12V +12V Si4497DY
J2 NC_01 NC_02 NC_03 /14V4 NC_04 NC_05 NC_06 GNDD NC_07 NC_08 Conn_01x10_Female
R3 Net-_D1-Pad2_ /14V4 10k
D1 /14V4 Net-_D1-Pad2_ 10V
U1 /14V4 Net-_D1-Pad2_ 15V
R8 Net-_Q3-Pad3_ Net-_D1-Pad2_ 10k
U3 +12V GNDD 15V
JP1 GNDD GND Jumper_2_Bridged
R6 Net-_Q2-Pad3_ Net-_Q3-Pad1_ 10k
J1 /14V4 Net-_J1-Pad2_ Conn_01x02_Female
D2 +12V Net-_D2-Pad2_ 1N4007
R7 Net-_J1-Pad2_ Net-_D2-Pad2_ 20
Q2 Net-_Q2-Pad1_ +12V Net-_Q2-Pad3_ BC807
R4 +12V Net-_Q2-Pad1_ 10k
Q1 Net-_Q1-Pad1_ GNDD Net-_Q1-Pad3_ BC817
R5 Net-_Q2-Pad1_ Net-_Q1-Pad3_ 4,7k
R2 Net-_Q1-Pad1_ GNDD 10k
R1 Net-_Q1-Pad1_ Net-_MCU_EN1-Pad1_ 1k
MCU_EN1 Net-_MCU_EN1-Pad1_ MCU_SUSTAIN
.end
